/* =========================================
* Top module wrapper of an accelerator role
*
* Author: Yisong Chang (changyisong@ict.ac.cn)
* Date: 29/01/2021
* Version: v0.0.1
*===========================================
*/

`timescale 10 ns / 1 ns

module role_top (
  input         aclk,
  input         aresetn,
  input		rtc_clock,

output [1:0]  m_axi_io_arid,
  output [30:0] m_axi_io_araddr,
  output [1:0]  m_axi_io_arburst,
  output [3:0]  m_axi_io_arcache,
  output [7:0]  m_axi_io_arlen,
  output [0:0]  m_axi_io_arlock,
  output [2:0]  m_axi_io_arprot,
  output [3:0]  m_axi_io_arqos,
  input         m_axi_io_arready,
  output [2:0] m_axi_io_arsize,
  output        m_axi_io_arvalid,
  output [1:0]  m_axi_io_awid,
  output [30:0] m_axi_io_awaddr,
  output [1:0] m_axi_io_awburst,
  output [3:0] m_axi_io_awcache,
  output [7:0] m_axi_io_awlen,
  output [0:0] m_axi_io_awlock,
  output [2:0] m_axi_io_awprot,
  output [3:0] m_axi_io_awqos,
  input         m_axi_io_awready,
  output [2:0] m_axi_io_awsize,
  output        m_axi_io_awvalid,
  input  [1:0]  m_axi_io_bid,
  output        m_axi_io_bready,
  input  [1:0]  m_axi_io_bresp,
  input         m_axi_io_bvalid,
  input  [1:0]  m_axi_io_rid,
  input  [63:0] m_axi_io_rdata,
  input         m_axi_io_rlast,
  output        m_axi_io_rready,
  input  [1:0]  m_axi_io_rresp,
  input         m_axi_io_rvalid,
  output [63:0] m_axi_io_wdata,
  output        m_axi_io_wlast,
  input         m_axi_io_wready,
  output [7:0]  m_axi_io_wstrb,
  output        m_axi_io_wvalid,
  
  
  output [35:0] m_axi_mem_araddr,
  output [1:0]  m_axi_mem_arburst,
  output [3:0]  m_axi_mem_arcache,
  output [7:0]  m_axi_mem_arlen,
  output [0:0]  m_axi_mem_arlock,
  output [2:0]  m_axi_mem_arprot,
  output [3:0]  m_axi_mem_arqos,
  input         m_axi_mem_arready,
  output [2:0]	m_axi_mem_arsize,
  output        m_axi_mem_arvalid,
  output [35:0]	m_axi_mem_awaddr,
  output [1:0]	m_axi_mem_awburst,
  output [3:0]	m_axi_mem_awcache,
  output [7:0]	m_axi_mem_awlen,
  output [0:0]	m_axi_mem_awlock,
  output [2:0]	m_axi_mem_awprot,
  output [3:0]	m_axi_mem_awqos,
  input         m_axi_mem_awready,
  output [2:0]	m_axi_mem_awsize,
  output        m_axi_mem_awvalid,
  output        m_axi_mem_bready,
  input  [1:0]  m_axi_mem_bresp,
  input         m_axi_mem_bvalid,
  input  [255:0] m_axi_mem_rdata,
  input         m_axi_mem_rlast,
  output        m_axi_mem_rready,
  input  [1:0]  m_axi_mem_rresp,
  input         m_axi_mem_rvalid,
  output [255:0] m_axi_mem_wdata,
  output        m_axi_mem_wlast,
  input         m_axi_mem_wready,
  output [31:0]  m_axi_mem_wstrb,
  output        m_axi_mem_wvalid,

  input  [19:0] s_axi_ctrl_araddr,
  input  [2:0]  s_axi_ctrl_arprot,
  output        s_axi_ctrl_arready,
  input         s_axi_ctrl_arvalid,
  input  [19:0] s_axi_ctrl_awaddr,
  input  [2:0]  s_axi_ctrl_awprot,
  output        s_axi_ctrl_awready,
  input         s_axi_ctrl_awvalid,
  input         s_axi_ctrl_bready,
  output [1:0]  s_axi_ctrl_bresp,
  output        s_axi_ctrl_bvalid,
  output [31:0] s_axi_ctrl_rdata,
  input         s_axi_ctrl_rready,
  output [1:0]  s_axi_ctrl_rresp,
  output        s_axi_ctrl_rvalid,
  input  [31:0] s_axi_ctrl_wdata,
  output        s_axi_ctrl_wready,
  input  [3:0]  s_axi_ctrl_wstrb,
  input         s_axi_ctrl_wvalid,

  input  [35:0] s_axi_dma_araddr,
  input  [13:0] s_axi_dma_arid,
  input  [1:0]  s_axi_dma_arburst,
  input  [3:0]  s_axi_dma_arcache,
  input  [7:0]  s_axi_dma_arlen,
  input  [0:0]  s_axi_dma_arlock,
  input  [2:0]  s_axi_dma_arprot,
  input  [3:0]  s_axi_dma_arqos,
  output        s_axi_dma_arready,
  input  [2:0]  s_axi_dma_arsize,
  input         s_axi_dma_arvalid,
  input  [35:0] s_axi_dma_awaddr,
  input  [13:0] s_axi_dma_awid,
  input  [1:0]  s_axi_dma_awburst,
  input  [3:0]  s_axi_dma_awcache,
  input  [7:0]  s_axi_dma_awlen,
  input  [0:0]  s_axi_dma_awlock,
  input  [2:0]  s_axi_dma_awprot,
  input  [3:0]  s_axi_dma_awqos,
  output        s_axi_dma_awready,
  input  [2:0]  s_axi_dma_awsize,
  input         s_axi_dma_awvalid,
  input         s_axi_dma_bready,
  output [1:0]  s_axi_dma_bresp,
  output        s_axi_dma_bvalid,
  output [13:0] s_axi_dma_bid,
  output [255:0]s_axi_dma_rdata,
  output        s_axi_dma_rlast,
  input         s_axi_dma_rready,
  output [1:0]  s_axi_dma_rresp,
  output        s_axi_dma_rvalid,
  output [13:0] s_axi_dma_rid,
  input  [255:0]s_axi_dma_wdata,
  input         s_axi_dma_wlast,
  output        s_axi_dma_wready,
  input  [31:0] s_axi_dma_wstrb,
  input         s_axi_dma_wvalid,

  output                m_axis_trace_tvalid,
  input                 m_axis_trace_tready,
  output  [512-1:0]     m_axis_trace_tdata,
  output  [512/8-1:0]   m_axis_trace_tkeep,
  output                m_axis_trace_tlast,

  input   [63:0]  s2r_intr
);

endmodule
