module xstop_wrapper (
  input          clk,
  input          rst,
  input          rtc_clk,

  output         dma_awready,
  input          dma_awvalid,
  input  [13:0]  dma_awid,
  input  [47:0]  dma_awaddr,
  input  [7:0]   dma_awlen,
  input  [2:0]   dma_awsize,
  input  [1:0]   dma_awburst,
  input          dma_awlock,
  input  [3:0]   dma_awcache,
  input  [2:0]   dma_awprot,
  input  [3:0]   dma_awqos,
  output         dma_wready,
  input          dma_wvalid,
  input  [255:0] dma_wdata,
  input  [31:0]  dma_wstrb,
  input          dma_wlast,
  input          dma_bready,
  output         dma_bvalid,
  output [13:0]  dma_bid,
  output [1:0]   dma_bresp,
  output         dma_arready,
  input          dma_arvalid,
  input  [13:0]  dma_arid,
  input  [47:0]  dma_araddr,
  input  [7:0]   dma_arlen,
  input  [2:0]   dma_arsize,
  input  [1:0]   dma_arburst,
  input          dma_arlock,
  input  [3:0]   dma_arcache,
  input  [2:0]   dma_arprot,
  input  [3:0]   dma_arqos,
  input          dma_rready,
  output         dma_rvalid,
  output [13:0]  dma_rid,
  output [255:0] dma_rdata,
  output [1:0]   dma_rresp,
  output         dma_rlast,
  input          peripheral_awready,
  output         peripheral_awvalid,
  output [1:0]   peripheral_awid,
  output [30:0]  peripheral_awaddr,
  output [7:0]   peripheral_awlen,
  output [2:0]   peripheral_awsize,
  output [1:0]   peripheral_awburst,
  output         peripheral_awlock,
  output [3:0]   peripheral_awcache,
  output [2:0]   peripheral_awprot,
  output [3:0]   peripheral_awqos,
  input          peripheral_wready,
  output         peripheral_wvalid,
  output [63:0]  peripheral_wdata,
  output [7:0]   peripheral_wstrb,
  output         peripheral_wlast,
  output         peripheral_bready,
  input          peripheral_bvalid,
  input  [1:0]   peripheral_bid,
  input  [1:0]   peripheral_bresp,
  input          peripheral_arready,
  output         peripheral_arvalid,
  output [1:0]   peripheral_arid,
  output [30:0]  peripheral_araddr,
  output [7:0]   peripheral_arlen,
  output [2:0]   peripheral_arsize,
  output [1:0]   peripheral_arburst,
  output         peripheral_arlock,
  output [3:0]   peripheral_arcache,
  output [2:0]   peripheral_arprot,
  output [3:0]   peripheral_arqos,
  output         peripheral_rready,
  input          peripheral_rvalid,
  input  [1:0]   peripheral_rid,
  input  [63:0]  peripheral_rdata,
  input  [1:0]   peripheral_rresp,
  input          peripheral_rlast,
  input          memory_awready,
  output         memory_awvalid,
  output [13:0]  memory_awid,
  output [47:0]  memory_awaddr,
  output [7:0]   memory_awlen,
  output [2:0]   memory_awsize,
  output [1:0]   memory_awburst,
  output         memory_awlock,
  output [3:0]   memory_awcache,
  output [2:0]   memory_awprot,
  output [3:0]   memory_awqos,
  input          memory_wready,
  output         memory_wvalid,
  output [255:0] memory_wdata,
  output [31:0]  memory_wstrb,
  output         memory_wlast,
  output         memory_bready,
  input          memory_bvalid,
  input  [13:0]  memory_bid,
  input  [1:0]   memory_bresp,
  input          memory_arready,
  output         memory_arvalid,
  output [13:0]  memory_arid,
  output [47:0]  memory_araddr,
  output [7:0]   memory_arlen,
  output [2:0]   memory_arsize,
  output [1:0]   memory_arburst,
  output         memory_arlock,
  output [3:0]   memory_arcache,
  output [2:0]   memory_arprot,
  output [3:0]   memory_arqos,
  output         memory_rready,
  input          memory_rvalid,
  input  [13:0]  memory_rid,
  input  [255:0] memory_rdata,
  input  [1:0]   memory_rresp,
  input          memory_rlast,

  output         riscv_halt,
  output         riscv_critical_error,
  output [63:0]  trace_cause,
  output [49:0]  trace_tval,
  output [2:0]   trace_priv,
  output [49:0]  trace_iaddr0,
  output [49:0]  trace_iaddr1,
  output [49:0]  trace_iaddr2,
  output [11:0]  trace_itype,
  output [20:0]  trace_iretire,
  output [2:0]   trace_ilastsize,

  input  [47:0]  rst_vec,
  input  [63:0]  ext_intrs
);
  wire [47:0] memory_araddr_raw;
  wire [47:0] memory_awaddr_raw;

  //assign memory_araddr = memory_araddr_raw - 48'h80000000;
  //assign memory_awaddr = memory_awaddr_raw - 48'h80000000;
  assign memory_araddr = memory_araddr_raw;
  assign memory_awaddr = memory_awaddr_raw;

  XSTop xstop(
    .io_clock(clk),
    .io_reset(rst),
    .io_rtc_clock(rtc_clk),
    .dma_awready(dma_awready),
    .dma_awvalid(dma_awvalid),
    .dma_awid(dma_awid),
    .dma_awaddr(dma_awaddr),
    .dma_awlen(dma_awlen),
    .dma_awsize(dma_awsize),
    .dma_awburst(dma_awburst),
    .dma_awlock(dma_awlock),
    .dma_awcache(dma_awcache),
    .dma_awprot(dma_awprot),
    .dma_awqos(dma_awqos),
    .dma_wready(dma_wready),
    .dma_wvalid(dma_wvalid),
    .dma_wdata(dma_wdata),
    .dma_wstrb(dma_wstrb),
    .dma_wlast(dma_wlast),
    .dma_bready(dma_bready),
    .dma_bvalid(dma_bvalid),
    .dma_bid(dma_bid),
    .dma_bresp(dma_bresp),
    .dma_arready(dma_arready),
    .dma_arvalid(dma_arvalid),
    .dma_arid(dma_arid),
    .dma_araddr(dma_araddr),
    .dma_arlen(dma_arlen),
    .dma_arsize(dma_arsize),
    .dma_arburst(dma_arburst),
    .dma_arlock(dma_arlock),
    .dma_arcache(dma_arcache),
    .dma_arprot(dma_arprot),
    .dma_arqos(dma_arqos),
    .dma_rready(dma_rready),
    .dma_rvalid(dma_rvalid),
    .dma_rid(dma_rid),
    .dma_rdata(dma_rdata),
    .dma_rresp(dma_rresp),
    .dma_rlast(dma_rlast),
    .peripheral_awready(peripheral_awready),
    .peripheral_awvalid(peripheral_awvalid),
    .peripheral_awid(peripheral_awid),
    .peripheral_awaddr(peripheral_awaddr),
    .peripheral_awlen(peripheral_awlen),
    .peripheral_awsize(peripheral_awsize),
    .peripheral_awburst(peripheral_awburst),
    .peripheral_awlock(peripheral_awlock),
    .peripheral_awcache(peripheral_awcache),
    .peripheral_awprot(peripheral_awprot),
    .peripheral_awqos(peripheral_awqos),
    .peripheral_wready(peripheral_wready),
    .peripheral_wvalid(peripheral_wvalid),
    .peripheral_wdata(peripheral_wdata),
    .peripheral_wstrb(peripheral_wstrb),
    .peripheral_wlast(peripheral_wlast),
    .peripheral_bready(peripheral_bready),
    .peripheral_bvalid(peripheral_bvalid),
    .peripheral_bid(peripheral_bid),
    .peripheral_bresp(peripheral_bresp),
    .peripheral_arready(peripheral_arready),
    .peripheral_arvalid(peripheral_arvalid),
    .peripheral_arid(peripheral_arid),
    .peripheral_araddr(peripheral_araddr),
    .peripheral_arlen(peripheral_arlen),
    .peripheral_arsize(peripheral_arsize),
    .peripheral_arburst(peripheral_arburst),
    .peripheral_arlock(peripheral_arlock),
    .peripheral_arcache(peripheral_arcache),
    .peripheral_arprot(peripheral_arprot),
    .peripheral_arqos(peripheral_arqos),
    .peripheral_rready(peripheral_rready),
    .peripheral_rvalid(peripheral_rvalid),
    .peripheral_rid(peripheral_rid),
    .peripheral_rdata(peripheral_rdata),
    .peripheral_rresp(peripheral_rresp),
    .peripheral_rlast(peripheral_rlast),
    .memory_awready(memory_awready),
    .memory_awvalid(memory_awvalid),
    .memory_awid(memory_awid),
    .memory_awaddr(memory_awaddr_raw),
    .memory_awlen(memory_awlen),
    .memory_awsize(memory_awsize),
    .memory_awburst(memory_awburst),
    .memory_awlock(memory_awlock),
    .memory_awcache(memory_awcache),
    .memory_awprot(memory_awprot),
    .memory_awqos(memory_awqos),
    .memory_wready(memory_wready),
    .memory_wvalid(memory_wvalid),
    .memory_wdata(memory_wdata),
    .memory_wstrb(memory_wstrb),
    .memory_wlast(memory_wlast),
    .memory_bready(memory_bready),
    .memory_bvalid(memory_bvalid),
    .memory_bid(memory_bid),
    .memory_bresp(memory_bresp),
    .memory_arready(memory_arready),
    .memory_arvalid(memory_arvalid),
    .memory_arid(memory_arid),
    .memory_araddr(memory_araddr_raw),
    .memory_arlen(memory_arlen),
    .memory_arsize(memory_arsize),
    .memory_arburst(memory_arburst),
    .memory_arlock(memory_arlock),
    .memory_arcache(memory_arcache),
    .memory_arprot(memory_arprot),
    .memory_arqos(memory_arqos),
    .memory_rready(memory_rready),
    .memory_rvalid(memory_rvalid),
    .memory_rid(memory_rid),
    .memory_rdata(memory_rdata),
    .memory_rresp(memory_rresp),
    .memory_rlast(memory_rlast),
    .nmi_0_0(0),
    .nmi_0_1(1),
    .io_sram_config(0),
    .io_pll0_lock(0),
    .io_pll0_ctrl_0(),
    .io_pll0_ctrl_1(),
    .io_pll0_ctrl_2(),
    .io_pll0_ctrl_3(),
    .io_pll0_ctrl_4(),
    .io_pll0_ctrl_5(),
    .io_systemjtag_jtag_TCK(0),
    .io_systemjtag_jtag_TMS(0),
    .io_systemjtag_jtag_TDI(0),
    .io_systemjtag_jtag_TDO_data(),
    .io_systemjtag_jtag_TDO_driven(),
    .io_systemjtag_reset(0),
    .io_systemjtag_mfr_id(0),
    .io_systemjtag_part_number(0),
    .io_systemjtag_version(0),
    .io_debug_reset(),
    .io_cacheable_check_req_0_valid(0),
    .io_cacheable_check_req_0_bits_addr(0),
    .io_cacheable_check_req_0_bits_size(0),
    .io_cacheable_check_req_0_bits_cmd(0),
    .io_cacheable_check_req_1_valid(0),
    .io_cacheable_check_req_1_bits_addr(0),
    .io_cacheable_check_req_1_bits_size(0),
    .io_cacheable_check_req_1_bits_cmd(0),
    .io_cacheable_check_resp_0_ld(),
    .io_cacheable_check_resp_0_st(),
    .io_cacheable_check_resp_0_instr(),
    .io_cacheable_check_resp_0_mmio(),
    .io_cacheable_check_resp_0_atomic(),
    .io_cacheable_check_resp_1_ld(),
    .io_cacheable_check_resp_1_st(),
    .io_cacheable_check_resp_1_instr(),
    .io_cacheable_check_resp_1_mmio(),
    .io_cacheable_check_resp_1_atomic(),
    .io_riscv_halt_0(riscv_halt),
    .io_riscv_critical_error_0(riscv_critical_error),
    .io_riscv_rst_vec_0(rst_vec),
    .io_traceCoreInterface_0_fromEncoder_enable(0),
    .io_traceCoreInterface_0_fromEncoder_stall(0),
    .io_traceCoreInterface_0_toEncoder_cause(trace_cause),
    .io_traceCoreInterface_0_toEncoder_tval(trace_tval),
    .io_traceCoreInterface_0_toEncoder_priv(trace_priv),
    .io_traceCoreInterface_0_toEncoder_iaddr({trace_iaddr2, trace_iaddr1, trace_iaddr0}),
    .io_traceCoreInterface_0_toEncoder_itype(trace_itype),
    .io_traceCoreInterface_0_toEncoder_iretire(trace_iretire),
    .io_traceCoreInterface_0_toEncoder_ilastsize(trace_ilastsize),
    .io_extIntrs(ext_intrs)
  );

endmodule
